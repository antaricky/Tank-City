module tank_yellow(output logic [4:0] rgb[0:127][0:15]);assign rgb = '{'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd11,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd10,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd9,4'd9,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd11,4'd11,4'd9,4'd9,4'd9,4'd11,4'd9,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd11,4'd9,4'd11,4'd11,4'd10,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd9,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd11,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd10,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd10,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd9,4'd9,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd11,4'd11,4'd9,4'd9,4'd9,4'd11,4'd9,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd9,4'd9,4'd9,4'd9,4'd11,4'd9,4'd11,4'd11,4'd10,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd9,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd11,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd9,4'd11,4'd9,4'd10,4'd10,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd9,4'd11,4'd10,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd10,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd10,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd9,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd9,4'd11,4'd9,4'd10,4'd10,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd9,4'd11,4'd10,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd10,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd11,4'd10,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd11,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd9,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd9,4'd9,4'd9,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd9,4'd11,4'd11,4'd10,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd11,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd10,4'd9,4'd11,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd9,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd9,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd9,4'd9,4'd9,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd9,4'd11,4'd11,4'd10,4'd11,4'd9,4'd9,4'd9,4'd9,4'd9,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd9,4'd11,4'd11,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd11,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd11,4'd10,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd11,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd11,4'd9,4'd11,4'd11,4'd11,4'd10,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd10,4'd10,4'd9,4'd10,4'd10,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd11,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd10,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd9,4'd9,4'd11,4'd11,4'd11,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd11,4'd9,4'd11,4'd11,4'd11,4'd10,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd11,4'd9,4'd11,4'd10,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd9,4'd11,4'd11,4'd10,4'd10,4'd11,4'd10,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd9,4'd9,4'd11,4'd11,4'd11,4'd11,4'd10,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd10,4'd10,4'd9,4'd0,4'd10,4'd10,4'd9,4'd10,4'd10,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd10,4'd11,4'd9,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd11,4'd11,4'd0,4'd0
},'{4'd0,4'd11,4'd10,4'd10,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd10,4'd10,4'd10,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd9,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
}};
endmodule
