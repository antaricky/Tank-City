module tank_silver(output logic [4:0] rgb[0:127][0:15]);assign rgb = '{'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd4,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd8,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd5,4'd5,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd5,4'd5,4'd5,4'd4,4'd5,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd4,4'd5,4'd4,4'd4,4'd8,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd4,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd8,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd8,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd5,4'd5,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd4,4'd4,4'd5,4'd5,4'd5,4'd4,4'd5,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd4,4'd5,4'd4,4'd4,4'd8,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd5,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd5,4'd4,4'd5,4'd8,4'd8,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd5,4'd4,4'd8,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd8,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd5,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd5,4'd4,4'd5,4'd8,4'd8,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd5,4'd4,4'd8,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd8,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd4,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd5,4'd5,4'd5,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd5,4'd4,4'd4,4'd8,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd8,4'd5,4'd4,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd5,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd5,4'd5,4'd5,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd5,4'd4,4'd4,4'd8,4'd4,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd4,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd4,4'd8,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd4,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd4,4'd5,4'd4,4'd4,4'd4,4'd8,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd8,4'd8,4'd5,4'd8,4'd8,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd4,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd8,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd5,4'd5,4'd4,4'd4,4'd4,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd4,4'd5,4'd4,4'd4,4'd4,4'd8,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd4,4'd5,4'd4,4'd8,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd5,4'd4,4'd4,4'd8,4'd8,4'd4,4'd8,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd5,4'd5,4'd4,4'd4,4'd4,4'd4,4'd8,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd8,4'd8,4'd5,4'd0,4'd8,4'd8,4'd5,4'd8,4'd8,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd8,4'd4,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd4,4'd4,4'd0,4'd0
},'{4'd0,4'd4,4'd8,4'd8,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd8,4'd8,4'd8,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
}};
endmodule
