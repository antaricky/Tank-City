module explosion(output logic [5:0] rgb[0:47][0:15]);
assign rgb = '{
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd16,5'd0,5'd15,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd16,5'd16,5'd15,5'd16,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd16,5'd15,5'd15,5'd0,5'd16,5'd15,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd15,5'd16,5'd15,5'd7,5'd15,5'd0,5'd7,5'd15,5'd15,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd16,5'd15,5'd7,5'd7,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd16,5'd7,5'd0,5'd7,5'd16,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd15,5'd15,5'd15,5'd7,5'd15,5'd7,5'd15,5'd15,5'd16,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd16,5'd16,5'd16,5'd16,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd0,5'd15,5'd16,5'd0,5'd16,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd16,5'd15,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd16,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd16,5'd0,5'd0,5'd15,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd16,5'd0,5'd15,5'd15,5'd16,5'd0,5'd0,5'd16,5'd15,5'd16,5'd0
},
'{
5'd0,5'd0,5'd16,5'd0,5'd15,5'd15,5'd16,5'd15,5'd16,5'd15,5'd15,5'd16,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd16,5'd7,5'd15,5'd15,5'd15,5'd15,5'd7,5'd15,5'd16,5'd16,5'd0,5'd0
},
'{
5'd0,5'd16,5'd15,5'd16,5'd16,5'd15,5'd7,5'd15,5'd0,5'd16,5'd15,5'd7,5'd15,5'd15,5'd15,5'd0
},
'{
5'd0,5'd0,5'd16,5'd15,5'd15,5'd15,5'd0,5'd7,5'd7,5'd7,5'd16,5'd15,5'd16,5'd16,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd7,5'd7,5'd7,5'd7,5'd0,5'd15,5'd16,5'd0,5'd16,5'd0
},
'{
5'd0,5'd0,5'd15,5'd15,5'd15,5'd16,5'd15,5'd7,5'd0,5'd7,5'd16,5'd15,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd15,5'd16,5'd16,5'd16,5'd7,5'd15,5'd0,5'd15,5'd15,5'd15,5'd7,5'd15,5'd15,5'd16,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd15,5'd15,5'd16,5'd16,5'd15,5'd16,5'd7,5'd16,5'd0,5'd0,5'd16,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd15,5'd16,5'd15,5'd16,5'd16,5'd15,5'd15,5'd16,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd16,5'd0,5'd16,5'd0,5'd15,5'd0,5'd16,5'd0,5'd0,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0
},
'{
5'd0,5'd15,5'd16,5'd0,5'd0,5'd15,5'd0,5'd15,5'd16,5'd0,5'd15,5'd0,5'd16,5'd15,5'd16,5'd0
},
'{
5'd0,5'd0,5'd16,5'd16,5'd0,5'd0,5'd16,5'd15,5'd16,5'd0,5'd16,5'd15,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd16,5'd16,5'd16,5'd15,5'd15,5'd16,5'd16,5'd16,5'd15,5'd16,5'd0,5'd0,5'd0
},
'{
5'd16,5'd0,5'd15,5'd15,5'd7,5'd15,5'd15,5'd0,5'd15,5'd16,5'd15,5'd15,5'd16,5'd0,5'd16,5'd0
},
'{
5'd0,5'd15,5'd0,5'd16,5'd15,5'd15,5'd7,5'd15,5'd15,5'd16,5'd15,5'd7,5'd15,5'd16,5'd0,5'd0
},
'{
5'd16,5'd0,5'd0,5'd16,5'd15,5'd7,5'd16,5'd7,5'd16,5'd0,5'd16,5'd15,5'd16,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd15,5'd15,5'd15,5'd7,5'd0,5'd7,5'd15,5'd15,5'd16,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd15,5'd15,5'd16,5'd15,5'd0,5'd7,5'd0,5'd0,5'd7,5'd0,5'd15,5'd15,5'd15,5'd15,5'd15
},
'{
5'd0,5'd0,5'd0,5'd16,5'd16,5'd15,5'd0,5'd7,5'd7,5'd0,5'd15,5'd16,5'd16,5'd16,5'd0,5'd0
},
'{
5'd0,5'd16,5'd0,5'd0,5'd15,5'd15,5'd7,5'd15,5'd15,5'd16,5'd7,5'd15,5'd16,5'd0,5'd0,5'd16
},
'{
5'd16,5'd0,5'd0,5'd15,5'd15,5'd7,5'd16,5'd15,5'd16,5'd16,5'd15,5'd15,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd0,5'd15,5'd15,5'd16,5'd16,5'd15,5'd15,5'd16,5'd15,5'd16,5'd0,5'd15,5'd16,5'd0,5'd0
},
'{
5'd0,5'd15,5'd16,5'd16,5'd16,5'd0,5'd16,5'd15,5'd16,5'd15,5'd16,5'd0,5'd0,5'd15,5'd16,5'd0
},
'{
5'd16,5'd16,5'd0,5'd0,5'd0,5'd0,5'd0,5'd15,5'd0,5'd0,5'd15,5'd0,5'd16,5'd0,5'd15,5'd16
},
'{
5'd0,5'd0,5'd0,5'd0,5'd16,5'd0,5'd0,5'd15,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
}};
endmodule
