module base(output logic [4:0] rgb[0:15][0:15]);assign rgb = '{'{4'd0,4'd1,4'd0,4'd1,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd2,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd2,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd1,4'd0,4'd0,4'd0,4'd1,4'd1,4'd2,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0
},'{4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd1,4'd2,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd0,4'd1,4'd0,4'd0,4'd1,4'd1,4'd2,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd1,4'd1,4'd2,4'd1,4'd1,4'd1,4'd0,4'd0,4'd1,4'd1,4'd0
},'{4'd0,4'd0,4'd0,4'd1,4'd1,4'd1,4'd2,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd1,4'd1,4'd1,4'd1,4'd1,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd1,4'd0,4'd1,4'd0,4'd1,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
}};
endmodule
