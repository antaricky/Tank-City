module steel(output logic [4:0] rgb[0:15][0:15]);assign rgb = '{'{4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4
},'{4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd1,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd4,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1
},'{4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1
},'{4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4
},'{4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd1,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd4,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1,4'd4,4'd4,4'd5,4'd5,4'd5,4'd5,4'd1,4'd1
},'{4'd4,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd4,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1
},'{4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd4,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1,4'd1
}};
endmodule
