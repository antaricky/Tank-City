module bullet(output logic [5:0] rgb[0:31][0:15]);
assign rgb = '{
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd4,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd4,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
}};
endmodule
