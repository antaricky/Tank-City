module tank_green(output logic [5:0] rgb[0:127][0:15]);
assign rgb = '{
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd14,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd12,5'd12,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd12,5'd12,5'd12,5'd14,5'd12,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd14,5'd12,5'd14,5'd14,5'd13,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd14,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd13,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd12,5'd12,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd14,5'd14,5'd12,5'd12,5'd12,5'd14,5'd12,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd12,5'd12,5'd12,5'd14,5'd12,5'd14,5'd14,5'd13,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd14,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd12,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd12,5'd14,5'd12,5'd13,5'd13,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd12,5'd14,5'd13,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd13,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd13,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd12,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd12,5'd14,5'd12,5'd13,5'd13,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd12,5'd14,5'd13,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd13,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd14,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd14,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd12,5'd12,5'd12,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd12,5'd14,5'd14,5'd13,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd13,5'd12,5'd14,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd12,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd12,5'd12,5'd12,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd12,5'd14,5'd14,5'd13,5'd14,5'd12,5'd12,5'd12,5'd12,5'd12,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd12,5'd14,5'd14,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd14,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd14,5'd13,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd14,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd14,5'd12,5'd14,5'd14,5'd14,5'd13,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd13,5'd13,5'd12,5'd13,5'd13,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd14,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd13,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd12,5'd12,5'd14,5'd14,5'd14,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd14,5'd12,5'd14,5'd14,5'd14,5'd13,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd14,5'd12,5'd14,5'd13,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd12,5'd14,5'd14,5'd13,5'd13,5'd14,5'd13,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd12,5'd12,5'd14,5'd14,5'd14,5'd14,5'd13,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd13,5'd13,5'd12,5'd0,5'd13,5'd13,5'd12,5'd13,5'd13,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd13,5'd14,5'd12,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd14,5'd14,5'd0,5'd0
},
'{
5'd0,5'd14,5'd13,5'd13,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd13,5'd13,5'd13,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd12,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
},
'{
5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0,5'd0
}};
endmodule
