module steel(output logic [5:0] rgb[0:15][0:15]);
assign rgb = '{
'{
5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4
},
'{
5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd1,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd4,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4
},
'{
5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd1,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd4,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1,5'd4,5'd4,5'd5,5'd5,5'd5,5'd5,5'd1,5'd1
},
'{
5'd4,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd4,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
},
'{
5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd4,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1,5'd1
}};
endmodule
