module palette(output logic [7:0] palette[0:15][0:2]);
assign palette = '{'{8'd0,8'd0,8'd1},'{8'd99,8'd99,8'd99},'{8'd107,8'd8,8'd0},'{8'd156,8'd74,8'd0},'{8'd173,8'd173,8'd173},'{8'd255,8'd255,8'd255},'{8'd90,8'd0,8'd123},'{8'd181,8'd49,8'd33},'{8'd0,8'd66,8'd74},'{8'd231,8'd231,8'd148},'{8'd107,8'd107,8'd0},'{8'd231,8'd156,8'd33},'{8'd181,8'd247,8'd206},'{8'd0,8'd82,8'd0},'{8'd0,8'd140,8'd49},'{8'd0,8'd0,8'd0}};
endmodule
