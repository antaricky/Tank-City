module tank_green(output logic [4:0] rgb[0:127][0:15]);assign rgb = '{'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd14,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd12,4'd12,4'd12,4'd12,4'd13,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd12,4'd12,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd14,4'd14,4'd12,4'd12,4'd12,4'd14,4'd12,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd12,4'd12,4'd12,4'd12,4'd14,4'd12,4'd14,4'd14,4'd13,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd12,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd12,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd14,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd13,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd12,4'd12,4'd12,4'd12,4'd13,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd12,4'd12,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd14,4'd14,4'd12,4'd12,4'd12,4'd14,4'd12,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd12,4'd12,4'd12,4'd12,4'd14,4'd12,4'd14,4'd14,4'd13,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd12,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd14,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd12,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd12,4'd14,4'd12,4'd13,4'd13,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd12,4'd14,4'd13,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd13,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd13,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd12,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd12,4'd14,4'd12,4'd13,4'd13,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd12,4'd14,4'd13,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd13,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd14,4'd13,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd14,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd12,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd12,4'd12,4'd12,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd12,4'd14,4'd14,4'd13,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd14,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd13,4'd12,4'd14,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd12,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd12,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd12,4'd12,4'd12,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd12,4'd14,4'd14,4'd13,4'd14,4'd12,4'd12,4'd12,4'd12,4'd12,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd12,4'd14,4'd14,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd14,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd14,4'd13,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd14,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd14,4'd12,4'd14,4'd14,4'd14,4'd13,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd13,4'd13,4'd12,4'd13,4'd13,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd14,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd13,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd12,4'd12,4'd14,4'd14,4'd14,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd14,4'd12,4'd14,4'd14,4'd14,4'd13,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd14,4'd12,4'd14,4'd13,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd12,4'd14,4'd14,4'd13,4'd13,4'd14,4'd13,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd12,4'd12,4'd14,4'd14,4'd14,4'd14,4'd13,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd13,4'd13,4'd12,4'd0,4'd13,4'd13,4'd12,4'd13,4'd13,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd13,4'd14,4'd12,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd14,4'd14,4'd0,4'd0
},'{4'd0,4'd14,4'd13,4'd13,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd13,4'd13,4'd13,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd12,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
}};
endmodule
