module tank_purple(output logic [4:0] rgb[0:127][0:15]);assign rgb = '{'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd7,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd6,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd5,4'd5,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd5,4'd5,4'd5,4'd7,4'd5,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd7,4'd5,4'd7,4'd7,4'd6,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd7,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd6,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd6,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd5,4'd5,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd7,4'd7,4'd5,4'd5,4'd5,4'd7,4'd5,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd5,4'd5,4'd5,4'd7,4'd5,4'd7,4'd7,4'd6,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd5,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd5,4'd7,4'd5,4'd6,4'd6,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd5,4'd7,4'd6,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd6,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd5,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd5,4'd7,4'd5,4'd6,4'd6,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd5,4'd7,4'd6,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd6,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd7,4'd6,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd5,4'd5,4'd5,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd5,4'd7,4'd7,4'd6,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd7,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd6,4'd5,4'd7,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd5,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd5,4'd5,4'd5,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd5,4'd7,4'd7,4'd6,4'd7,4'd5,4'd5,4'd5,4'd5,4'd5,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd5,4'd7,4'd7,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd7,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd7,4'd6,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd7,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd7,4'd5,4'd7,4'd7,4'd7,4'd6,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd6,4'd6,4'd5,4'd6,4'd6,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd7,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd6,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd5,4'd5,4'd7,4'd7,4'd7,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd7,4'd5,4'd7,4'd7,4'd7,4'd6,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd7,4'd5,4'd7,4'd6,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd5,4'd7,4'd7,4'd6,4'd6,4'd7,4'd6,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd5,4'd5,4'd7,4'd7,4'd7,4'd7,4'd6,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd6,4'd6,4'd5,4'd0,4'd6,4'd6,4'd5,4'd6,4'd6,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd6,4'd7,4'd5,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd7,4'd7,4'd0,4'd0
},'{4'd0,4'd7,4'd6,4'd6,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd6,4'd6,4'd6,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd5,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
},'{4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0,4'd0
}};
endmodule
